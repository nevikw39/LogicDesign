module PAT(clk, reset, data, flag);
	
	input clk, reset, data;
	output flag;
	
endmodule
