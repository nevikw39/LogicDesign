`timescale 1ns / 1ps
`define SDFFILE "build/ALU.sdf"

module tb();

	parameter n = 16;
	parameter m = 4;
	parameter delay = 4;

	reg [n - 1: 0] A, B;
	reg Cin;
	reg [m - 1: 0] Mode;
	
	wire [n - 1: 0] Y;
	wire Cout, Overflow;

	reg [n - 1: 0] Y_correct;
	reg Cout_correct, Overflow_correct;

	ALU alu(A, B, Cin, Mode, Y, Cout, Overflow);

	initial begin
		`ifdef SDF
			$sdf_annotate(`SDFFILE, alu);
		`endif
	end

	integer file, r, i;
	reg [n - 1: 0] score;
	wire special_Mode;
	assign special_Mode = Mode == 4'b0100 || Mode == 4'b0101;

	initial begin
		file = $fopen("./data.txt", "r");
		score = 16'd0;
		i = 0;
		while (!$feof(file)) begin
			#delay;
			r = $fscanf(file, "%b %b %b %b %b %b %b", A, B, Cin, Mode, Y_correct, Cout_correct, Overflow_correct);
			#delay;
			if (Y === Y_correct && (!special_Mode || (special_Mode && Cout == Cout_correct && Overflow == Overflow_correct))) begin
				score = score + 16'd1;
			end
			else begin
				$display("WA: Testcase %2d", i);
				$display("A: (%b, %d), B: (%b, %d), Cin: %b, Mode: %d, ", A, $signed(A), B, $signed(B), Cin, Mode);
				$display("Your output,    Y: (%b, %d), Cout: %b, Overflow: %b", Y, $signed(Y), special_Mode ? Cout : 1'bx, special_Mode ? Overflow : 1'bx);
				$display("Correct output, Y: (%b, %d), Cout: %b, Overflow: %b", Y_correct, $signed(Y_correct), special_Mode ? Cout_correct : 1'bx, special_Mode ? Overflow_correct : 1'bx);
				$display("-----------------------------------");
			end
			i = i + 1;
		end
		#delay;
		$display("Total score: %d / %d", score, 64);
		if (score == 64) begin
			$display("AC");
		end
	end

endmodule
